module vsql

// ISO/IEC 9075-2:2016(E), 14.8, <delete statement: positioned>
//
// Delete a row of a table.
