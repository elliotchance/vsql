// ISO/IEC 9075-2:2016(E), 6.9, <set function specification>

module vsql

// Format
//~
//~ <set function specification> /* Expr */ ::=
//~     <aggregate function>
