// ISO/IEC 9075-2:2016(E), 6.28, <value expression>

module vsql

// Format
//~
//~ <value expression> /* Expr */ ::=
//~     <common value expression>
//~   | <boolean value expression>
//~
//~ <common value expression> /* Expr */ ::=
//~     <numeric value expression>
//~   | <string value expression>
//~   | <datetime value expression>
