// ISO/IEC 9075-2:2016(E), 8.1, <predicate>

module vsql

// Format
//~
//~ <predicate> /* Expr */ ::=
//~     <comparison predicate>
//~   | <between predicate>
//~   | <like predicate>
//~   | <similar predicate>
//~   | <null predicate>
