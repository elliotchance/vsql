module vsql

// ISO/IEC 9075-2:2016(E), 7.2, <row value expression>
//
// Specify a row value.
