// ISO/IEC 9075-2:2016(E), 6.35, <datetime value expression>

module vsql

// Format
//~
//~ <datetime value expression> /* Expr */ ::=
//~     <datetime term>
//~
//~ <datetime term> /* Expr */ ::=
//~     <datetime factor>
//~
//~ <datetime factor> /* Expr */ ::=
//~     <datetime primary>
//~
//~ <datetime primary> /* Expr */ ::=
//~     <value expression primary>
//~   | <datetime value function>
