module vsql

// ISO/IEC 9075-2:2016(E), 7.5, <from clause>
//
// Specify a table derived from one or more tables.
