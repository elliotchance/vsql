// ISO/IEC 9075-2:2016(E), 8.21, <search condition>

module vsql

// Format
//~
//~ <search condition> /* Expr */ ::=
//~     <boolean value expression>
