module vsql

fn is_reserved_word(word string) bool {
	reserved_words := ['ABS', 'ACOS', 'ALL', 'ALLOCATE', 'ALTER', 'AND', 'ANY', 'ARE', 'ARRAY',
		'ARRAY_AGG', 'ARRAY_MAX_CARDINALITY', 'AS', 'ASENSITIVE', 'ASIN', 'ASYMMETRIC', 'AT', 'ATAN',
		'ATOMIC', 'AUTHORIZATION', 'AVG', 'BEGIN', 'BEGIN_FRAME', 'BEGIN_PARTITION', 'BETWEEN',
		'BIGINT', 'BINARY', 'BLOB', 'BOOLEAN', 'BOTH', 'BY', 'CALL', 'CALLED', 'CARDINALITY',
		'CASCADED', 'CASE', 'CAST', 'CEIL', 'CEILING', 'CHAR', 'CHAR_LENGTH', 'CHARACTER',
		'CHARACTER_LENGTH', 'CHECK', 'CLASSIFIER', 'CLOB', 'CLOSE', 'COALESCE', 'COLLATE', 'COLLECT',
		'COLUMN', 'COMMIT', 'CONDITION', 'CONNECT', 'CONSTRAINT', 'CONTAINS', 'CONVERT', 'COPY',
		'CORR', 'CORRESPONDING', 'COS', 'COSH', 'COUNT', 'COVAR_POP', 'COVAR_SAMP', 'CREATE', 'CROSS',
		'CUBE', 'CUME_DIST', 'CURRENT', 'CURRENT_CATALOG', 'CURRENT_DATE',
		'CURRENT_DEFAULT_TRANSFORM_GROUP', 'CURRENT_PATH', 'CURRENT_ROLE', 'CURRENT_ROW',
		'CURRENT_SCHEMA', 'CURRENT_TIME', 'CURRENT_TIMESTAMP', 'CURRENT_PATH', 'CURRENT_ROLE',
		'CURRENT_TRANSFORM_GROUP_FOR_TYPE', 'CURRENT_USER', 'CURSOR', 'CYCLE', 'DATE', 'DAY',
		'DEALLOCATE', 'DEC', 'DECIMAL', 'DECFLOAT', 'DECLARE', 'DEFAULT', 'DEFINE', 'DELETE',
		'DENSE_RANK', 'DEREF', 'DESCRIBE', 'DETERMINISTIC', 'DISCONNECT', 'DISTINCT', 'DOUBLE',
		'DROP', 'DYNAMIC', 'EACH', 'ELEMENT', 'ELSE', 'EMPTY', 'END', 'END_FRAME', 'END_PARTITION',
		'END-EXEC', 'EQUALS', 'ESCAPE', 'EVERY', 'EXCEPT', 'EXEC', 'EXECUTE', 'EXISTS', 'EXP',
		'EXTERNAL', 'EXTRACT', 'FALSE', 'FETCH', 'FILTER', 'FIRST_VALUE', 'FLOAT', 'FLOOR', 'FOR',
		'FOREIGN', 'FRAME_ROW', 'FREE', 'FROM', 'FULL', 'FUNCTION', 'FUSION', 'GET', 'GLOBAL',
		'GRANT', 'GROUP', 'GROUPING', 'GROUPS', 'HAVING', 'HOLD', 'HOUR', 'IDENTITY', 'IN',
		'INDICATOR', 'INITIAL', 'INNER', 'INOUT', 'INSENSITIVE', 'INSERT', 'INT', 'INTEGER',
		'INTERSECT', 'INTERSECTION', 'INTERVAL', 'INTO', 'IS', 'JOIN', 'JSON_ARRAY', 'JSON_ARRAYAGG',
		'JSON_EXISTS', 'JSON_OBJECT', 'JSON_OBJECTAGG', 'JSON_QUERY', 'JSON_TABLE',
		'JSON_TABLE_PRIMITIVE', 'JSON_VALUE', 'LAG', 'LANGUAGE', 'LARGE', 'LAST_VALUE', 'LATERAL',
		'LEAD', 'LEADING', 'LEFT', 'LIKE', 'LIKE_REGEX', 'LISTAGG', 'LN', 'LOCAL', 'LOCALTIME',
		'LOCALTIMESTAMP', 'LOG', 'LOG10', 'LOWER', 'MATCH', 'MATCH_NUMBER', 'MATCH_RECOGNIZE',
		'MATCHES', 'MAX', 'MEMBER', 'MERGE', 'METHOD', 'MIN', 'MINUTE', 'MOD', 'MODIFIES', 'MODULE',
		'MONTH', 'MULTISET', 'NATIONAL', 'NATURAL', 'NCHAR', 'NCLOB', 'NEW', 'NO', 'NONE',
		'NORMALIZE', 'NOT', 'NTH_VALUE', 'NTILE', 'NULL', 'NULLIF', 'NUMERIC', 'OCTET_LENGTH',
		'OCCURRENCES_REGEX', 'OF', 'OFFSET', 'OLD', 'OMIT', 'ON', 'ONE', 'ONLY', 'OPEN', 'OR',
		'ORDER', 'OUT', 'OUTER', 'OVER', 'OVERLAPS', 'OVERLAY', 'PARAMETER', 'PARTITION', 'PATTERN',
		'PER', 'PERCENT', 'PERCENT_RANK', 'PERCENTILE_CONT', 'PERCENTILE_DISC', 'PERIOD', 'PORTION',
		'POSITION', 'POSITION_REGEX', 'POWER', 'PRECEDES', 'PRECISION', 'PREPARE', 'PRIMARY',
		'PROCEDURE', 'PTF', 'RANGE', 'RANK', 'READS', 'REAL', 'RECURSIVE', 'REF', 'REFERENCES',
		'REFERENCING', 'REGR_AVGX', 'REGR_AVGY', 'REGR_COUNT', 'REGR_INTERCEPT', 'REGR_R2',
		'REGR_SLOPE', 'REGR_SXX', 'REGR_SXY', 'REGR_SYY', 'RELEASE', 'RESULT', 'RETURN', 'RETURNS',
		'REVOKE', 'RIGHT', 'ROLLBACK', 'ROLLUP', 'ROW', 'ROW_NUMBER', 'ROWS', 'RUNNING', 'SAVEPOINT',
		'SCOPE', 'SCROLL', 'SEARCH', 'SECOND', 'SEEK', 'SELECT', 'SENSITIVE', 'SESSION_USER', 'SET',
		'SHOW', 'SIMILAR', 'SIN', 'SINH', 'SKIP', 'SMALLINT', 'SOME', 'SPECIFIC', 'SPECIFICTYPE',
		'SQL', 'SQLEXCEPTION', 'SQLSTATE', 'SQLWARNING', 'SQRT', 'START', 'STATIC', 'STDDEV_POP',
		'STDDEV_SAMP', 'SUBMULTISET', 'SUBSET', 'SUBSTRING', 'SUBSTRING_REGEX', 'SUCCEEDS', 'SUM',
		'SYMMETRIC', 'SYSTEM', 'SYSTEM_TIME', 'SYSTEM_USER', 'TABLE', 'TABLESAMPLE', 'TAN', 'TANH',
		'THEN', 'TIME', 'TIMESTAMP', 'TIMEZONE_HOUR', 'TIMEZONE_MINUTE', 'TO', 'TRAILING',
		'TRANSLATE', 'TRANSLATE_REGEX', 'TRANSLATION', 'TREAT', 'TRIGGER', 'TRIM', 'TRIM_ARRAY',
		'TRUE', 'TRUNCATE', 'UESCAPE', 'UNION', 'UNIQUE', 'UNKNOWN', 'UNNEST', 'UPDATE', 'UPPER',
		'USER', 'USING', 'VALUE', 'VALUES', 'VALUE_OF', 'VAR_POP', 'VAR_SAMP', 'VARBINARY', 'VARCHAR',
		'VARYING', 'VERSIONING', 'WHEN', 'WHENEVER', 'WHERE', 'WIDTH_BUCKET', 'WINDOW', 'WITH',
		'WITHIN', 'WITHOUT', 'YEAR']

	return word.to_upper() in reserved_words
}

fn is_non_reserved_word(word string) bool {
	non_reserved_words := ['A', 'ABSOLUTE', 'ACTION', 'ADA', 'ADD', 'ADMIN', 'AFTER', 'ALWAYS',
		'ASC', 'ASSERTION', 'ASSIGNMENT', 'ATTRIBUTE', 'ATTRIBUTES', 'BEFORE', 'BERNOULLI', 'BREADTH',
		'C', 'CASCADE', 'CATALOG', 'CATALOG_NAME', 'CHAIN', 'CHAINING', 'CHARACTER_SET_CATALOG',
		'CHARACTER_SET_NAME', 'CHARACTER_SET_SCHEMA', 'CHARACTERISTICS', 'CHARACTERS', 'CLASS_ORIGIN',
		'COBOL', 'COLLATION', 'COLLATION_CATALOG', 'COLLATION_NAME', 'COLLATION_SCHEMA', 'COLUMNS',
		'COLUMN_NAME', 'COMMAND_FUNCTION', 'COMMAND_FUNCTION_CODE', 'COMMITTED', 'CONDITIONAL',
		'CONDITION_NUMBER', 'CONNECTION', 'CONNECTION_NAME', 'CONSTRAINT_CATALOG', 'CONSTRAINT_NAME',
		'CONSTRAINT_SCHEMA', 'CONSTRAINTS', 'CONSTRUCTOR', 'CONTINUE', 'CURSOR_NAME', 'DATA',
		'DATETIME_INTERVAL_CODE', 'DATETIME_INTERVAL_PRECISION', 'DEFAULTS', 'DEFERRABLE', 'DEFERRED',
		'DEFINED', 'DEFINER', 'DEGREE', 'DEPTH', 'DERIVED', 'DESC', 'DESCRIBE_CATALOG',
		'DESCRIBE_NAME', 'DESCRIBE_PROCEDURE_SPECIFIC_CATALOG', 'DESCRIBE_PROCEDURE_SPECIFIC_NAME',
		'DESCRIBE_PROCEDURE_SPECIFIC_SCHEMA', 'DESCRIBE_SCHEMA', 'DESCRIPTOR', 'DIAGNOSTICS',
		'DISPATCH', 'DOMAIN', 'DYNAMIC_FUNCTION', 'DYNAMIC_FUNCTION_CODE', 'ENCODING', 'ENFORCED',
		'ERROR', 'EXCLUDE', 'EXCLUDING', 'EXPRESSION', 'FINAL', 'FINISH', 'FINISH_CATALOG',
		'FINISH_NAME', 'FINISH_PROCEDURE_SPECIFIC_CATALOG', 'FINISH_PROCEDURE_SPECIFIC_NAME',
		'FINISH_PROCEDURE_SPECIFIC_SCHEMA', 'FINISH_SCHEMA', 'FIRST', 'FLAG', 'FOLLOWING', 'FORMAT',
		'FORTRAN', 'FOUND', 'FULFILL', 'FULFILL_CATALOG', 'FULFILL_NAME',
		'FULFILL_PROCEDURE_SPECIFIC_CATALOG', 'FULFILL_PROCEDURE_SPECIFIC_NAME',
		'FULFILL_PROCEDURE_SPECIFIC_SCHEMA', 'FULFILL_SCHEMA', 'G', 'GENERAL', 'GENERATED', 'GO',
		'GOTO', 'GRANTED', 'HAS_PASS_THROUGH_COLUMNS', 'HAS_PASS_THRU_COLS', 'HIERARCHY', 'IGNORE',
		'IMMEDIATE', 'IMMEDIATELY', 'IMPLEMENTATION', 'INCLUDING', 'INCREMENT', 'INITIALLY', 'INPUT',
		'INSTANCE', 'INSTANTIABLE', 'INSTEAD', 'INVOKER', 'ISOLATION', 'IS_PRUNABLE', 'JSON', 'K',
		'KEEP', 'KEY', 'KEYS', 'KEY_MEMBER', 'KEY_TYPE', 'LAST', 'LENGTH', 'LEVEL', 'LOCATOR',
		'M', 'MAP', 'MATCHED', 'MAXVALUE', 'MESSAGE_LENGTH', 'MESSAGE_OCTET_LENGTH', 'MESSAGE_TEXT',
		'MINVALUE', 'MORE', 'MUMPS', 'NAME', 'NAMES', 'NESTED', 'NESTING', 'NEXT', 'NFC', 'NFD',
		'NFKC', 'NFKD', 'NORMALIZED', 'NULLABLE', 'NULLS', 'NUMBER', 'OBJECT', 'OCTETS', 'OPTION',
		'OPTIONS', 'ORDERING', 'ORDINALITY', 'OTHERS', 'OUTPUT', 'OVERFLOW', 'OVERRIDING', 'P',
		'PAD', 'PARAMETER_MODE', 'PARAMETER_NAME', 'PARAMETER_ORDINAL_POSITION',
		'PARAMETER_SPECIFIC_CATALOG', 'PARAMETER_SPECIFIC_NAME', 'PARAMETER_SPECIFIC_SCHEMA',
		'PARTIAL', 'PASCAL', 'PASS', 'PASSING', 'PAST', 'PATH', 'PLACING', 'PLAN', 'PLI', 'PRECEDING',
		'PRESERVE', 'PRIOR', 'PRIVATE', 'PRIVATE_PARAMETERS', 'PRIVATE_PARAMS_S', 'PRIVILEGES',
		'PRUNE', 'PUBLIC', 'QUOTES', 'READ', 'RELATIVE', 'REPEATABLE', 'RESPECT', 'RESTART',
		'RESTRICT', 'RETURNED_CARDINALITY', 'RETURNED_LENGTH', 'RETURNED_OCTET_LENGTH',
		'RETURNED_SQLSTATE', 'RETURNING', 'RETURNS_ONLY_PASS_THROUGH', 'RET_ONLY_PASS_THRU', 'ROLE',
		'ROUTINE', 'ROUTINE_CATALOG', 'ROUTINE_NAME', 'ROUTINE_SCHEMA', 'ROW_COUNT', 'SCALAR',
		'SCALE', 'SCHEMA', 'SCHEMA_NAME', 'SCOPE_CATALOG', 'SCOPE_NAME', 'SCOPE_SCHEMA', 'SECTION',
		'SECURITY', 'SELF', 'SEQUENCE', 'SERIALIZABLE', 'SERVER_NAME', 'SESSION', 'SETS', 'SIMPLE',
		'SIZE', 'SOURCE', 'SPACE', 'SPECIFIC_NAME', 'START_CATALOG', 'START_NAME',
		'START_PROCEDURE_SPECIFIC_CATALOG', 'START_PROCEDURE_SPECIFIC_NAME',
		'START_PROCEDURE_SPECIFIC_SCHEMA', 'START_SCHEMA', 'STATE', 'STATEMENT', 'STRING',
		'STRUCTURE', 'STYLE', 'SUBCLASS_ORIGIN', 'T', 'TABLE_NAME', 'TABLE_SEMANTICS', 'TEMPORARY',
		'THROUGH', 'TIES', 'TOP_LEVEL_COUNT', 'TRANSACTION', 'TRANSACTION_ACTIVE',
		'TRANSACTIONS_COMMITTED', 'TRANSACTIONS_ROLLED_BACK', 'TRANSFORM', 'TRANSFORMS',
		'TRIGGER_CATALOG', 'TRIGGER_NAME', 'TRIGGER_SCHEMA', 'TYPE', 'UNBOUNDED', 'UNCOMMITTED',
		'UNCONDITIONAL', 'UNDER', 'UNNAMED', 'USAGE', 'USER_DEFINED_TYPE_CATALOG',
		'USER_DEFINED_TYPE_CODE', 'USER_DEFINED_TYPE_NAME', 'USER_DEFINED_TYPE_SCHEMA', 'UTF16',
		'UTF32', 'UTF8', 'VIEW', 'WORK', 'WRAPPER', 'WRITE', 'ZONE']

	return word.to_upper() in non_reserved_words
}

fn is_key_word(word string) bool {
	return is_reserved_word(word) || is_non_reserved_word(word)
}
