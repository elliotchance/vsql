// ISO/IEC 9075-2:2016(E), 7.12, <where clause>

module vsql

// Format
//~
//~ <where clause> /* Expr */ ::=
//~     WHERE <search condition>   -> expr
