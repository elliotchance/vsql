module vsql

// ISO/IEC 9075-2:2016(E), 5.1, <SQL terminal character>
//
// # Function
//
// Define the terminal symbols of the SQL language and the elements of strings.
//
// # Format
//~
//~ <left paren> ::= "("
//~
//~ <right paren> ::= ")"
//~
//~ <asterisk> /* string */ ::=
//~   "*"
//~
//~ <plus sign> /* string */ ::=
//~   "+"
//~
//~ <comma> ::= ","
//~
//~ <minus sign> /* string */ ::=
//~   "-"
//~
//~ <period> ::= "."
//~
//~ <solidus> /* string */ ::=
//~   "/"
//~
//~ <colon> ::=
//~   ":"
//~
//~ <less than operator> ::= "<"
//~
//~ <equals operator> ::= "="
//~
//~ <greater than operator> ::= ">"
