module vsql

// ISO/IEC 9075-2:2016(E), 6.9, <set function specification>
//
// # Function
//
// Specify a value derived by the application of a function to an argument.
//
// # Format
//~
//~ <set function specification> /* AggregateFunction */ ::=
//~     <aggregate function>
