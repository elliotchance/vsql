// ISO/IEC 9075-2:2016(E), 14.3, <cursor specification>

module vsql

// Format
//~
//~ <cursor specification> /* Stmt */ ::=
//~     <query expression>   -> Stmt
