// ISO/IEC 9075-2:2016(E), 7.2, <row value expression>

module vsql

// Format
//~
//~ <table row value expression> /* Expr */ ::=
//~     <row value constructor>
//~
//~ <contextually typed row value expression> /* []Expr */ ::=
//~   <contextually typed row value constructor>
//~
//~ <row value predicand> /* Expr */ ::=
//~   <row value constructor predicand>
