// ISO/IEC 9075-2:2016(E), 11.6, <table constraint definition>

module vsql

// Format
//~
//~ <table constraint definition> /* TableElement */ ::=
//~   <table constraint>
//~
//~ <table constraint> /* TableElement */ ::=
//~   <unique constraint definition>
