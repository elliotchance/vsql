// ISO/IEC 9075-2:2016(E), 5.1, <SQL terminal character>

module vsql

// Format
//~
//~ <left paren> ::= "("
//~
//~ <right paren> ::= ")"
//~
//~ <asterisk> /* string */ ::=
//~   "*"
//~
//~ <plus sign> /* string */ ::=
//~   "+"
//~
//~ <comma> ::= ","
//~
//~ <minus sign> /* string */ ::=
//~   "-"
//~
//~ <period> ::= "."
//~
//~ <solidus> /* string */ ::=
//~   "/"
//~
//~ <colon> ::=
//~   ":"
//~
//~ <less than operator> ::= "<"
//~
//~ <equals operator> ::= "="
//~
//~ <greater than operator> ::= ">"
