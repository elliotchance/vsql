module vsql

// ISO/IEC 9075-2:2016(E), 20.7, <prepare statement>
//
// Prepare a statement for execution.
