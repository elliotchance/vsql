module vsql

// ISO/IEC 9075-2:2016(E), 7.2, <row value expression>
//
// # Function
//
// Specify a row value.
//
// # Format
//~
//~ <table row value expression> /* RowValueConstructor */ ::=
//~     <row value constructor>
//~
//~ <contextually typed row value expression> /* ContextuallyTypedRowValueConstructor */ ::=
//~   <contextually typed row value constructor>
//~
//~ <row value predicand> /* RowValueConstructorPredicand */ ::=
//~   <row value constructor predicand>
