module main

import vsql

fn main() {
	vsql.main_()
}
