// ISO/IEC 9075-2:2016(E), 14.8, <delete statement: positioned>

module vsql

// Format
//~
//~ <target table> /* Identifier */ ::=
//~     <table name>
