module vsql

// ISO/IEC 9075-2:2016(E), 14.3, <cursor specification>
//
// # Function
//
// Define a result set.
//
// # Format
//~
//~ <cursor specification> /* Stmt */ ::=
//~     <query expression>   -> Stmt
